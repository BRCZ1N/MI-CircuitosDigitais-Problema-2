module modulo_status_dig_2(d,clock,clr,prst,q)

	input d,clock,clr,prst;
	output q;

endmodule 