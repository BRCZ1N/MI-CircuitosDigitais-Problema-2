module modulo_contador_mod_6(t,clk,clr,q);

	input t,clk,clr;
	output reg q;
	

endmodule 