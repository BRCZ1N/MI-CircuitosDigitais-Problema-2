module modulo_contador_2bits(d,clock,clr,prst,q)

	input d,clock,clr,prst;
	output q;

endmodule 