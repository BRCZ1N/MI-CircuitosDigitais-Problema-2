module modulo_demux1_16(d,clock,clr,prst,q)

	input d,clock,clr,prst;
	output q;

endmodule 