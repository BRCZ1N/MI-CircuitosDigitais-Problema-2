module modulo_demux4_1(d,clock,clr,prst,q)

	input d,clock,clr,prst;
	output q;

endmodule 