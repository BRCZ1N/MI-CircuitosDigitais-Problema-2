module modulo_seletor_reg(d,clock,clr,prst,q);

	input d,clock,clr,prst;
	output q;

endmodule 