module modulo_demux16_1(d,clock,clr,prst,q)

	input d,clock,clr,prst;
	output q;

endmodule 