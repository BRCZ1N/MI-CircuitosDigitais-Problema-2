module modulo_decodificador_bcd_ex_7Seg(d,clock,clr,prst,q);

	input d,clock,clr,prst;
	output q;

endmodule 