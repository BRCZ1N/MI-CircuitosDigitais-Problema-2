module modulo_decodificador_bcd_ex_7seg_ac(d,clock,clr,prst,q);

	input d,clock,clr,prst;
	output q;

endmodule 