module pbl(d,clock,clr,prst,q);

	input d,clock,clr,prst;
	output q;

endmodule 