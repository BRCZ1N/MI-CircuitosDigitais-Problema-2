module modulo_coord_coluna(d,clock,clr,prst,q)

	input d,clock,clr,prst;
	output q;

endmodule 